library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity banco_de_regs is
    port(
        read_reg1   : in unsigned(15 downto 0);
        read_reg2   : in unsigned(15 downto 0);
        value       : in unsigned(15 downto 0);
        write_reg   : in unsigned(15 downto 0);
        write_en    : in std_logic;
        clk         : in std_logic;
        rst         : in std_logic;
        read_data1  : out unsigned(15 downto 0);
        read_data2  : out unsigned(15 downto 0)
    );
end entity;

architecture a_banco_de_regs of banco_de_regs is

    component reg16bits
        port(
            clk         : in std_logic;
            rst         : in std_logic;
            wr_en       : in std_logic;
            data_in     : in  unsigned(15 downto 0);
            data_out    : out unsigned(15 downto 0)
        );
    end component;

    constant reg0           : unsigned(15 downto 0) := "0000000000000000";
    constant reg1           : unsigned(15 downto 0) := "0000000000000001";
    constant reg2           : unsigned(15 downto 0) := "0000000000000010";
    constant reg3           : unsigned(15 downto 0) := "0000000000000011";
    constant reg4           : unsigned(15 downto 0) := "0000000000000100";
    constant reg5           : unsigned(15 downto 0) := "0000000000000101";
    constant reg6           : unsigned(15 downto 0) := "0000000000000110";
    constant reg7           : unsigned(15 downto 0) := "0000000000000111";
    constant error_value    : unsigned(15 downto 0) := "1111111111111111";
    constant zero           : unsigned(15 downto 0) := "0000000000000000"

    -- Single clock, reset and only write in 1 register per time
    signal clk_s, rst_s     : std_logic;    
    signal data_in_s        : unsigned(15 downto 0);

    -- Register 0
    signal wr_en_0_s        : std_logic;
    signal data_out_0_s     : unsigned(15 downto 0);

    -- Register 1
    signal wr_en_1_s        : std_logic;
    signal data_out_1_s     : unsigned(15 downto 0);

    -- Register 2
    signal wr_en_2_s        : std_logic;
    signal data_out_2_s     : unsigned(15 downto 0);

    -- Register 3
    signal wr_en_3_s        : std_logic;
    signal data_out_3_s     : unsigned(15 downto 0);

    -- Register 4
    signal wr_en_4_s        : std_logic;
    signal data_out_4_s     : unsigned(15 downto 0);

    -- Register 5
    signal wr_en_5_s        : std_logic;
    signal data_out_5_s     : unsigned(15 downto 0);

    -- Register 6
    signal wr_en_6_s        : std_logic;
    signal data_out_6_s     : unsigned(15 downto 0);

    -- Register 7
    signal wr_en_7_s        : std_logic;
    signal data_out_7_s     : unsigned(15 downto 0);

begin
    register_0 : reg16bits
    port map(
        clk         => clk_s,
        rst         => rst_s,
        wr_en       => wr_en_0_s,
        data_in     => data_in_s,
        data_out    => data_out_0_s,
    );

    register_1 : reg16bits
    port map(
        clk         => clk_s,
        rst         => rst_s,
        wr_en       => wr_en_1_s,
        data_in     => data_in_s,
        data_out    => data_out_1_s,
    );

    register_2 : reg16bits
    port map(
        clk         => clk_s,
        rst         => rst_s,
        wr_en       => wr_en_2_s,
        data_in     => data_in_s,
        data_out    => data_out_2_s,
    );

    register_3 : reg16bits
    port map(
        clk         => clk_s,
        rst         => rst_s,
        wr_en       => wr_en_3_s,
        data_in     => data_in_s,
        data_out    => data_out_3_s,
    );

    register_4 : reg16bits
    port map(
        clk         => clk_s,
        rst         => rst_s,
        wr_en       => wr_en_4_s,
        data_in     => data_in_s,
        data_out    => data_out_4_s,
    );

    register_5 : reg16bits
    port map(
        clk         => clk_s,
        rst         => rst_s,
        wr_en       => wr_en_5_s,
        data_in     => data_in_s,
        data_out    => data_out_5_s,
    );

    register_6 : reg16bits
    port map(
        clk         => clk_s,
        rst         => rst_s,
        wr_en       => wr_en_6_s,
        data_in     => data_in_s,
        data_out    => data_out_6_s,
    );

    register_7 : reg16bits
    port map(
        clk         => clk_s,
        rst         => rst_s,
        wr_en       => wr_en_7_s,
        data_in     => data_in_s,
        data_out    => data_out_7_s,
    );

    read_data1_p : process(clk, rst)
    begin
        if read_reg1 = reg0 then                    -- Case register 0
            read_data1 <= data_out_0_s;
        elsif read_reg1 = reg1 then                 -- Case register 1
            read_data1 <= data_out_1_s;
        elsif read_reg1 = reg2 then                 -- Case register 2
            read_data1 <= data_out_2_s;
        elsif read_reg1 = reg3 then                 -- Case register 3
            read_data1 <= data_out_3_s;
        elsif read_reg1 = reg4 then                 -- Case register 4
            read_data1 <= data_out_4_s;
        elsif read_reg1 = reg5 then                 -- Case register 5
            read_data1 <= data_out_5_s;
        elsif read_reg1 = reg6 then                 -- Case register 6
            read_data1 <= data_out_6_s;
        elsif read_reg1 = reg7 then                 -- Case register 7
            read_data1 <= data_out_7_s;
        else
            read_data1 <= error_value;
        end if;
    end process read_data1_p;

    read_data2_p : process(clk, rst)
    begin
        if read_reg2 = reg0 then                    -- Case register 0
            read_data2 <= data_out_0_s;
        elsif read_reg2 = reg1 then                 -- Case register 1
            read_data2 <= data_out_1_s;
        elsif read_reg2 = reg2 then                 -- Case register 2
            read_data2 <= data_out_2_s;
        elsif read_reg2 = reg3 then                 -- Case register 3
            read_data2 <= data_out_3_s;
        elsif read_reg2 = reg4 then                 -- Case register 4
            read_data2 <= data_out_4_s;
        elsif read_reg2 = reg5 then                 -- Case register 5
            read_data2 <= data_out_5_s;
        elsif read_reg2 = reg6 then                 -- Case register 6
            read_data2 <= data_out_6_s;
        elsif read_reg2 = reg7 then                 -- Case register 7
            read_data2 <= data_out_7_s;
        else
            read_data2 <= error_value;
        end if;
    end process read_data2_p;

end architecture